//========================================================================
// Basic.v
//========================================================================
// A basic in-order, single-issue decoder that implements TinyRV1

`ifndef HW_DECODE_DECODE_VARIANTS_BASIC_V
`define HW_DECODE_DECODE_VARIANTS_BASIC_V

`include "defs/ISA.v"
`include "intf/F__DIntf.v"

module Decode #(
  parameter p_addr_bits = 32,
  parameter p_inst_bits = 32
)(
  input  logic clk,
  input  logic rst,

  //----------------------------------------------------------------------
  // F <-> D Interface
  //----------------------------------------------------------------------

  F__DIntf.D_intf F,

  //----------------------------------------------------------------------
  // D <-> X Interface
  //----------------------------------------------------------------------

  D__XIntf.D_intf Ex
);

  //----------------------------------------------------------------------
  // Pipeline registers for F interface
  //----------------------------------------------------------------------

  typedef struct packed {
    logic                   val;
    logic [p_inst_bits-1:0] inst;
    logic [p_addr_bits-1:0] pc;
  } F_input;

  F_input F_reg;
  F_input F_reg_next
  logic   F_xfer;

  always_ff @( posedge clk ) begin
    if ( rst )
      F_reg <= '{ val: 1'b0, inst: 'x, pc: 'x };
    else
      F_reg <= F_reg_next;
  end

  always_comb begin
    F_xfer = F.val & F.rdy;

    if ( F_xfer )
      F_reg_next = '{ val: 1'b1, inst: F.inst, pc: F.pc };
    else
      F_reg_next = '{ val: 1'b0, inst: 'x, pc: 'x };
  end



endmodule

`endif // HW_DECODE_DECODE_VARIANTS_BASIC_V
